package types ;
  
typedef struct {
int pid ;
} packet ;

endpackage : types 
// create package types here

